/*
:name: behavior_of_randomization_methods_0
:description: static random variables test
:tags: 18.6.3
*/

class a;
    static rand int b;
    constraint c { b > 5; b < 12; }
endclass

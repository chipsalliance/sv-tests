/*
:name: empty_test_2
:description: Test
:tags: 5.3 5.4
*/
			
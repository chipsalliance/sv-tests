/*
:name: class_test_25
:description: Test
:tags: 6.15 8.3
*/
package Package;
	interface class Bar; endclass
endpackage

class Foo implements Package::Bar; endclass

module test;
endmodule

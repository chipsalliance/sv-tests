/*
:name: class_member_test_14
:description: Test
:tags: 8.3
*/
class myclass;
function integer subroutine;
  input a;
  subroutine = a+42;
endfunction
endclass

module test;
endmodule

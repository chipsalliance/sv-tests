/*
:name: typedef_test_23
:description: Test
:tags: 6.18
*/
typedef bit[3:0] num_t;
typedef enum num_t {
  Global = 4'h2,
  Local = 4'h3
} myenum_fwd;

module test;
endmodule

/*
:name: 22.4--include_basic
:description: Test
:tags: 22.4
:type: preprocessing parsing
*/
`include "dummy_include.sv"
module top ();
endmodule

/*
:name: class_member_test_29
:description: Test
:should_fail: 1
:tags: 8.3
*/
class myclass;
function void shifter;
  for (int shft_idx  = 0 ; shft_idx < n_bits ) begin
  end
endfunction
endclass

/*
:name: typedef_test_22
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef enum uvec8_t;
typedef enum {
  Global = 2,
  Local = 3
} uvec8_t;

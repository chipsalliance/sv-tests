/*
:name: typedef_test_15
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef struct packed {
  [4:0] some_member;
} mystruct_t;
/*
:name: uvm_files
:description: basic UVM test
:tags: uvm
:timeout: 100
*/


/*
:name: class_test_39
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class macros_as_class_item;
 `moobar(,)
 `zoobar(  ,  )
 `zootar(12,)
 `zoojar(,34)
endclass
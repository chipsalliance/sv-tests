/*
:name: vector_vectored
:description: vectored vector tests
:should_fail: 0
:tags: 6.9.2
*/
module top();
	logic vectored [15:0] a;

	a = 12;
endmodule

/*
:name: typedef_test_24
:description: Test
:tags: 6.18
*/
typedef struct {
  int sample;
  int tile;
} tuple_t;

module test;
endmodule

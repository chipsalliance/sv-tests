/*
:name: preproc_test_2
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`include "preproc_test_2.svh"
`ifndef SUCCESS
Didn't successfully include preproc_test_2.svh!
`endif
`ifndef SANITY
`define SANITY
`endif

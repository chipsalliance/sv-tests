/*
:name: class_member_test_25
:description: Test
:tags: 8.3
*/
class myclass;
extern virtual function integer subroutine;
endclass

function integer myclass::subroutine; endfunction

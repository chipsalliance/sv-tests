// -*- coding: utf-8 -*-
//
// Copyright (C) 2020 The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
// SPDX-License-Identifier: ISC

package testbench_pkg;
   `include "uvm_macros.svh"
   import uvm_pkg::*;
   
//   import testbench_agent_pkg::*;

//   `include "testbench_env_config.svh"
//   `include "testbench_env.svh"
//   `include "custom_report_server.svh"
//   `include "testbench_base_test.svh"
//   `include "cto_scoreboard_config.svh"
//   `include "cto_scoreboard.svh"
     `include "cto_monitor.svh"
endpackage

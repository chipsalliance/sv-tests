/*
:name: constraint_blocks_0
:description: constraint blocks test
:tags: 18.5
*/

class a;
    rand int b;
    constraint c { b == 0; }
endclass

/*
:name: class_member_test_3
:description: Test
:tags: 8.3
*/
class myclass;
extern task subtask(int arg);
endclass

task myclass::subtask(int arg); endtask

module test;
endmodule

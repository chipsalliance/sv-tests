/*
:name: class_test_6
:description: Test
:tags: 6.15 8.3
*/
class Bar; endclass
class Foo extends Bar; endclass

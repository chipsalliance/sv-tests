/*
:name: localparam
:description: localparam without type specifier
:tags: 6.20.4
*/
module top();
	localparam p = 123;
endmodule

/*
:name: typedef_test_3
:description: Test
:tags: 6.18
*/
typedef reg[1:0] quartet[1:0];

module test;
endmodule

/*
:name: preproc_test_7
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`define INCEPTION(a, b, c) \
  (a*b-c)

module test;
endmodule

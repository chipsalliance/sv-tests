/*
:name: typedef_test_1
:description: Test
:tags: 6.18
*/
typedef reg[3:0] quartet;

module test;
endmodule

/*
:name: typedef_test_0
:description: Test
:tags: 6.18
*/
typedef i_am_a_type_really;

typedef int i_am_a_type_really;

// Multiple forward typedefs are allowed.
typedef i_am_a_type_really;
typedef i_am_a_type_really;

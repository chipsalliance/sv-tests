/*
:name: rand_modifier
:description: rand modifier test
:tags: 18.4.1
*/

class a;
    rand int b;
endclass

// -*- coding: utf-8 -*-
//
// Copyright (C) 2020 The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
// SPDX-License-Identifier: ISC


package test_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"

   import sys_uvc_pkg::*;
   import axi_agent_pkg::*;
   import axi_env_pkg::*;
   import axi_seq_pkg::*;
   import common_pkg::*;

   `include "axi_test_list.svh"
endpackage

/*
:name: struct_test_0
:description: Test
:tags: 7.2
*/
typedef struct mystruct_fwd;

typedef struct { logic a; logic b; } mystruct_fwd;
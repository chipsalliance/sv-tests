/*
:name: number_test_6
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
module test;
parameter integer foo = 1'b0;
endmodule

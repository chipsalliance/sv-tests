// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: attributes-operator
:description: Assing attributes to an operator
:tags: 5.12
*/

module top();
  logic [7:0] a;
  logic [7:0] b;
  logic [7:0] c;

  initial begin
    a = b + (* mode = "cla" *) c;
  end

endmodule

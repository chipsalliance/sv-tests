// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: localparam_type_decl
:description: Declare a type with a localparam
:tags: 6.23
*/
module top ;

localparam type testtype = logic;

testtype t;

endmodule

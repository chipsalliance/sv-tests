/*
:name: number_test_7
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 1'B0;

module test;
endmodule

/*
:name: number_test_19
:description: Test
:should_fail: 0
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 16'b`DIGITS(bar);
/*
:name: number_test_47
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 32 'o 7;

module test;
endmodule

/*
:name: set_membership_0
:description: set membership test
:tags: 18.5.3
*/

class a;
    rand int b;
    constraint c { b inside {3, 10}; }
endclass

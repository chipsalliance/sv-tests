/*
:name: typedef_test_19
:description: Test
:tags: 6.18
*/
typedef enum {
  Global = 2,
  Local = 3
} myenum_fwd;
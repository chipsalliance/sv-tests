// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: preproc_test_2
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`include "preproc_test_2.svh"
`ifndef SUCCESS
"Didn't successfully include preproc_test_2.svh!"
`endif
`ifndef SANITY
`define SANITY
`endif

module test;
endmodule

/*
:name: class_member_test_8
:description: Test
:tags: 8.3
*/
class myclass;
extern protected virtual task subtask(int arg);
endclass

task myclass::subtask(int arg);
endtask

/*
:name: iface_class_test_0
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic;
endclass

module test;
endmodule

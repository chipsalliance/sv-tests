/*
:name: class_member_test_6
:description: Test
:tags: 8.3
*/
class myclass;
extern protected task subtask(int arg);
endclass

task myclass::subtask(int arg); endtask
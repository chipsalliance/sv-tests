/*
:name: class_member_test_18
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subroutine(input bit x);
endclass

function void myclass::subroutine(input bit x);
endfunction

/*
:name: class_member_test_7
:description: Test
:tags: 8.3
*/
class myclass;
extern virtual protected task subtask(int arg);
endclass

task myclass::subtask(int arg);
endtask

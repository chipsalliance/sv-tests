/*
:name: typedef_test_7
:description: Test
:tags: 6.18
*/
typedef struct { int i, j, k; bit b, c, d; } mystruct;

module test;
endmodule

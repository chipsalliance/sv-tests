/*
:name: class_test_4
:description: Test
:tags: 6.15 8.3
*/
virtual class Foo; endclass

module test;
endmodule

/*
:name: pure_constraint_1
:description: pure constraint test
:tags: 18.5.2 uvm
*/

import uvm_pkg::*;
`include "uvm_macros.svh"

virtual class a;
    pure constraint c;
endclass

class a2 extends a;
    rand int b2;
    constraint c { b2 == 5; }
endclass

class env extends uvm_env;

  a2 obj = new;

  function new(string name, uvm_component parent = null);
    super.new(name, parent);
  endfunction
  
  task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    begin
      obj.randomize();
      if(obj.b2 == 5) begin
        `uvm_info("RESULT", $sformatf("b2 = %0d SUCCESS", obj.b2), UVM_LOW);
      end else begin
        `uvm_info("RESULT", $sformatf("b2 = %0d FAILED", obj.b2), UVM_LOW);
      end
    end
    phase.drop_objection(this);
  endtask: run_phase
  
endclass

module top;

  env environment;

  initial begin
    environment = new("env");
    run_test();
  end
  
endmodule

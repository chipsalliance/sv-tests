/*
:name: class_member_test_41
:description: Test
:tags: 8.3
*/
class constructible;
function new ();
endfunction : new
endclass

module test;
endmodule

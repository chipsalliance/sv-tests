/*
:name: class_test_38
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class macros_as_class_item;
 `moobar()
 `zoobar(  )
 `zootar(
)
endclass
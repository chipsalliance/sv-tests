/*
:name: 22.11--pragma-invalid
:description: Test
:should_fail_because: The pragma specification is identified by the pragma_name, which follows the `pragma directive.
:tags: 22.11
:type: preprocessing
*/
`pragma

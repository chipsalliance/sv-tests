/*
:name: class_member_test_15
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subroutine;
endclass

function void myclass::subroutine;
endfunction

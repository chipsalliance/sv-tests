/*
:name: 22.12--line-illegal-5
:description: Missing filename 
:should_fail_because: Missing filename 
:tags: 22.12
:type: preprocessing
*/
`line 1

/*
:name: localparam_int
:description: localparam integer type
:tags: 6.20.4
*/
module top();
	localparam int p = 123;
endmodule

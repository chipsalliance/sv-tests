/*
:name: class_member_test_0
:description: Test
:tags: 8.3
*/
class myclass;
task subtask;
endtask
endclass

module test;
endmodule

/*
:name: localparam_uint
:description: localparam unsigned typed
:tags: 6.20.4
*/
module top();
	localparam int unsigned q = 123;
endmodule

/*
:name: class_member_test_3
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern task automatic subtask(arg_type arg);
endclass
/*
:name: 22.9--unconnected_drive-invalid-1
:description: Test
:should_fail_because: The directive `unconnected_drive takes one of two arguments - pull1 or pull0.
:tags: 22.9
:type: simulation
*/
`unconnected_drive
`nounconnected_drive

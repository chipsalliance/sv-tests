// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: ferror_function
:description: $ferror test
:tags: 21.3
:type: simulation elaboration parsing
*/
module top();

initial begin
	int fd;
	string str;
	integer errno;
	fd = $fopen("tmp.txt", "w");
	errno = $ferror(fd, str);
	$display(errno);
	$display(str);
	$fclose(fd);
end

endmodule

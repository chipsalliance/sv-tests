/*
:name: class_test_58
:description: Test
:tags: 6.15 8.3
*/
typedef int data_type_or_module_type;

class fields_with_modifiers;
  const static data_type_or_module_type foo1 = 4'hf;
  static const data_type_or_module_type foo3 = 1, foo4 = 2;
endclass

module test;
endmodule

/*
:name: static_constraint_blocks_0
:description: static constraint blocks test
:tags: 18.5.11
*/

class a;
    rand int b;

    static constraint c1 { b == 5; }
endclass



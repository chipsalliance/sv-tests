/*
:name: class_test_55
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Driver;
  Packet pNP [*];
  Packet pNP1 [*];
  Packet pNP2 [*];
  Packet pNP3 [*];
endclass

/*
:name: number_test_8
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 1 'b 0;

module test;
endmodule

/*
:name: class_member_test_22
:description: Test
:should_fail: 1
:tags: 8.3
*/
class myclass;
extern function sometype #(N+1)[N:0]subr(ducktype #(3) x);
endclass

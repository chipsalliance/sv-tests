/*
:name: empty_test_1
:description: Test
:tags: 5.3 5.4
*/
    
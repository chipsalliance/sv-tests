/*
:name: number_test_14
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 4'bzzzz;

module test;
endmodule

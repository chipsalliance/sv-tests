// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: class_member_test_40
:description: Test
:tags: 8.3
:unsynthesizable: 1
*/
class constructible;
function new ();
endfunction
endclass

module test;
endmodule

/*
:name: number_test_0
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter foo = 0;

module test;
endmodule

/*
:name: number_test_23
:description: Test
:should_fail: 0
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = `WIDTH'b`DIGITS;
/*
:name: number_test_43
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 'o 0;

module test;
endmodule

/*
:name: class_test_60
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
`ifdef DEBUGGER
`ifdef VERBOSE
`endif
`endif
endclass

module test;
endmodule

/*
:name: typedef_test_18
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef struct {
  rand bit i;
  randc integer b[k:0];
} randstruct;

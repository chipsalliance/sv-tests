// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: finish_task
:description: $finish test
:tags: 20.2
:unsynthesizable: 1
*/
module top();

initial
	$finish;

endmodule

/*
:name: unconnected-drive
:description: Unconnected drive keywords
:tags: 5.6.4
:type: preprocessing
*/


`unconnected_drive pull1

module ts();
endmodule

`nounconnected_drive

/*
:name: class_test_11
:description: Test
:tags: 6.15 8.3
*/
class Foo #(int N, int P);
endclass

module test;
endmodule

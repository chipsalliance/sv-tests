/*
:name: class_member_test_39
:description: Test
:tags: 8.3
*/
class constructible;
function new;
endfunction
endclass

module test;
endmodule

/*
:name: union_test_0
:description: Test
:tags: 7.3
*/
typedef union myunion_fwd;

typedef union { logic a; logic b; } myunion_fwd;

/*
:name: class_test_15
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo #(type KeyType=int, Int=int);
endclass
/*
:name: iface_class_test_6
:description: Test
:should_fail: 0
:tags: 8.3 8.26
*/
interface class base_ic;
typedef int[3:0] quartet;
typedef string string_type;
endclass
/*
:name: class_test_55
:description: Test
:tags: 6.15 8.3
*/
class Packet;
endclass

class Driver;
  Packet pNP [*];
  Packet pNP1 [* ];
  Packet pNP2 [ *];
  Packet pNP3 [ * ];
endclass

// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: one_net_assign
:description: simple net declaration assignment test
:tags: 10.3.1
:type: simulation elaboration parsing
*/
module top(input a, output b);

assign b = a;

endmodule

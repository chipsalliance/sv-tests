/*
:name: empty_test_0
:description: Test
:tags: 5.3 5.4
*/

/*
:name: typedef_test_19
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef enum {
  Global = 2,
  Local = 3
} myenum_fwd;
/*
:name: empty_test_5
:description: Test
:tags: 5.3 5.4
*/
/* comment */

/*
:name: number_test_27
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 32'D1;

module test;
endmodule

/*
:name: unconnected-drive
:description: Unconnected drive keywords
:should_fail: 0
:tags: 5.6.4
*/

`nounconnected_drive
`unconnected_drive

module ts();
endmodule

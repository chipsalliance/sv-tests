/*
:name: iface_class_test_1
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic;
endclass : base_ic

module test;
endmodule

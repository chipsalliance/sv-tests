/*
:name: class_test_48
:description: Test
:tags: 6.15 8.3
*/
class pp_as_class_item;
 `undef EVIL_MACRO
endclass

module test;
endmodule

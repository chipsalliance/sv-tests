/*
:name: class_member_test_4
:description: Test
:tags: 8.3
*/
class myclass;
extern virtual task subtask(int arg);
endclass

task myclass::subtask(int arg); endtask

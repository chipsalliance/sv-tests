/*
:name: class_test_1
:description: Test
:tags: 6.15 8.3
*/
class Foo; endclass

module test;
endmodule

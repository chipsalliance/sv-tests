/*
:name: empty_test_4
:description: Test
:tags: 5.3 5.4
*/
// comment

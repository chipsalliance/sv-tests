/*
:name: compiler_directives_preprocessor_macro_0
:description: Read preprocessing macro from template (:defines: marker)
:tags: 5.6.4
:defines: TEST_VAR
*/

`ifdef TEST_VAR
`else
TEST_VAR parsed not correctly from template
`endif

// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: shortreal
:description: shortreal type tests
:tags: 6.12
:unsynthesizable: 1
*/
module top();
	shortreal a = 0.5;
endmodule

/*
:name: typedef_test_21
:description: Test
:tags: 6.18
*/
typedef enum bit[3:0] {
  Global = 4'h2,
  Local = 4'h3
} myenum_fwd;

module test;
endmodule

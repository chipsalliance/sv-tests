/*
:name: randc_modifier
:description: randc modifier test
:tags: 18.4.2
*/

class a;
    randc int b;
endclass

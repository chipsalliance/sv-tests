/*
:name: basic
:description: Test dynamic arrays support
:should_fail: 0
:tags: 7.5
*/
module top ();

bit [7:0] arr[];

endmodule

/*
:name: number_test_68
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 32'Sh7;

module test;
endmodule

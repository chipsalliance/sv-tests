/*
:name: class_test_57
:description: Test
:tags: 6.15 8.3
*/
typedef int data_type_or_module_type;

class fields_with_modifiers;
  const data_type_or_module_type foo1 = 4'hf;
  static data_type_or_module_type foo3, foo4;
endclass

module test;
endmodule

/*
:name: string_itoa
:description: string.itoa()  tests
:should_fail: 0
:tags: 6.16.11
*/
module top();
	string a;
	a.itoa(12);
endmodule

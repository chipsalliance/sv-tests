/*
:name: class_test_9
:description: Test
:tags: 6.15 8.3
*/
class Foo #(int N);
endclass

module test;
endmodule

/*
:name: typedef_test_4
:description: Test
:tags: 6.18
*/
typedef enum { RED, GREEN, BLUE } colors;

module test;
endmodule

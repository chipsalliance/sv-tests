/*
:name: class_test_69
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
  int num_packets;
`ifdef DEBUGGER
`elsif BORED
`else
  string source_name;
  string dest_name;
`endif
  int router_size;
endclass

module test;
endmodule

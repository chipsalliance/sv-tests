/*
:name: typedef_test_8
:description: Test
:tags: 6.18
*/
typedef bit some_other_type;
typedef some_other_type myalias;

module test;
endmodule

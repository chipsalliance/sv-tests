/*
:name: class_test_0
:description: Test
:tags: 6.15 8.3
*/
class semicolon_classy; ; ;;; ; ; ;endclass

module test;
endmodule

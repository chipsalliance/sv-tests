/*
:name: class_test_28
:description: Test
:tags: 6.15 8.3
*/

class Base; endclass
interface class Bar; endclass

class Foo extends Base implements Bar; endclass

module test;
endmodule

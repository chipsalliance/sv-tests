/*
:name: class_member_test_16
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function automatic void subroutine;
endclass
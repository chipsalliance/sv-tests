/*
:name: typedef_test_22
:description: Test
:tags: 6.18
*/
typedef enum uvec8_t;
typedef enum {
  Global = 2,
  Local = 3
} uvec8_t;

/*
:name: class_test_35
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class zzxx;
extern function /*automatic*/ void set_port(int ap);
endclass

/*
:name: class_member_test_18
:description: Test
:tags: 8.3
*/
class myclass;
typedef logic bool;
extern function void subroutine(input bool x);
endclass

function void myclass::subroutine(input bool x); endfunction

module test;
endmodule

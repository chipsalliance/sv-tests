/*
:name: class_test_7
:description: Test
:tags: 6.15 8.3
*/
package Package;
  class Bar; endclass
endpackage

class Foo extends Package::Bar; endclass
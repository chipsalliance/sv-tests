// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: class_test_55
:description: Test
:tags: 6.15 8.3
:unsynthesizable: 1
*/
class Packet;
endclass

class Driver;
  Packet pNP [*];
  Packet pNP1 [* ];
  Packet pNP2 [ *];
  Packet pNP3 [ * ];
endclass

module test;
endmodule

/*
:name: typedef_test_10
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef data_t my_array_t [*];

// -*- coding: utf-8 -*-
//
// Copyright (C) 2020 The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
// SPDX-License-Identifier: ISC

`ifndef _AXI_SEQ_LIST_SVH_
`define _AXI_SEQ_LIST_SVH_

`include "axi_base_seq.svh"
`include "axi_wrap_seq.svh"
`include "tb_axi_seq.svh"

`endif

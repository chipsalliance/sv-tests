/*
:name: basic
:description: Test memories support
:should_fail: 0
:tags: 7.4.4
*/
module top ();

// one-dimensinal array with elements of types
// reg, logic, bit
logic [7:0] mem [0:255];

endmodule

/*
:name: typedef_test_5
:description: Test
:tags: 6.18
*/
typedef union { int i; bit b; } bint;

module test;
endmodule

/*
:name: class_test_18
:description: Test
:tags: 6.15 8.3
*/
class Foo #(type IFType=virtual interface x_if);
endclass

module test;
endmodule

// -*- coding: utf-8 -*-
//
// Copyright (C) 2020 The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
// SPDX-License-Identifier: ISC

package testbench_pkg;
   `include "uvm_macros.svh"
   import uvm_pkg::*;

     `include "cto_monitor.svh"
endpackage

/*
:name: one_net_assign
:description: simple net declaration assignment test
:tags: 10.3.1
:type: parsing simulation
*/
module top(input a, output b);

assign b = a;

endmodule

/*
:name: class_member_test_9
:description: Test
:tags: 8.3
*/
class myclass;
typedef int arg_type;
extern local static task subtask(arg_type arg);
endclass

task myclass::subtask(arg_type arg); endtask

module test;
endmodule

/*
:name: localparam_string
:description: localparam string typed
:tags: 6.20.4
*/
module top();
	localparam s1 = "foo";
	localparam string s2 = "bar";
endmodule

/*
:name: typedef_test_8__bad
:description: Test
:should_fail_because: defining a type using an undefined type
:tags: 6.18
:type: simulation
*/
// some_other_type is not defined
typedef some_other_type myalias;

module test;
endmodule

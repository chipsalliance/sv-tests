// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: static_constraint_blocks_0
:description: static constraint blocks test
:tags: 18.5.11
:unsynthesizable: 1
*/

class a;
    rand int b;

    static constraint c1 { b == 5; }
endclass

/*
:name: empty_test_3
:description: Test
:tags: 5.3 5.4
*/



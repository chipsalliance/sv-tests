/*
:name: 22.9--unconnected_drive-invalid-3
:description: Test
:should_fail_because: use a strength keyword with `nounconnected_drive macro
:tags: 22.9
:type: simulation
*/
`unconnected_drive pull0 
`nounconnected_drive pull0

/*
:name: 22.12--line-illegal-4
:description: The level parameter shall be 0, 1, or 2
:should_fail_because: The level parameter shall be 0, 1, or 2
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile"
